module dmem(
    addr,
    dataW,
    clk,
    dataB,
    MemRW,
);

    input [31:0] addr;
    input [31:0] dataW;
    input clk;
    input MemRW;
    output reg [31:0] dataB;

    parameter read = 0;
    parameter write = 1;

    reg [31:0] mem_arr [0:31];
    
	initial begin
	    mem_arr[0]=32'b00000000000000000000000000000000;
		mem_arr[1]=32'b00000000000000000000000000000000;
		mem_arr[2]=32'b00000000000000000000000000000000;
		mem_arr[3]=32'b00000000000000000000000000000000;
		mem_arr[4]=32'b00000000000000000000000000000000;
		mem_arr[5]=32'b00000000000000000000000000000000;
		mem_arr[6]=32'b00000000000000000000000000000000;
		mem_arr[7]=32'b00000000000000000000000000000000;
		mem_arr[8]=32'b00000000000000000000000000000000;
		mem_arr[9]=32'b00000000000000000000000000000000;
		mem_arr[10]=32'b00000000000000000000000000000000;
		mem_arr[11]=32'b00000000000000000000000000000000;
		mem_arr[12]=32'b00000000000000000000000000000000;
		mem_arr[13]=32'b00000000000000000000000000000000;
		mem_arr[14]=32'b00000000000000000000000000000000;
		mem_arr[15]=32'b00000000000000000000000000000000;
		mem_arr[16]=32'b00000000000000000000000000000000;
		mem_arr[17]=32'b00000000000000000000000000000000;
		mem_arr[18]=32'b00000000000000000000000000000000;
		mem_arr[19]=32'b00000000000000000000000000000000;
		mem_arr[20]=32'b00000000000000000000000000000000;
		mem_arr[21]=32'b00000000000000000000000000000000;
		mem_arr[22]=32'b00000000000000000000000000000000;
		mem_arr[23]=32'b00000000000000000000000000000000;
		mem_arr[25]=32'b00000000000000000000000000000000;
		mem_arr[26]=32'b00000000000000000000000000000000;
		mem_arr[27]=32'b00000000000000000000000000000000;
		mem_arr[28]=32'b00000000000000000000000000000000;
		mem_arr[29]=32'b00000000000000000000000000000000;
		mem_arr[30]=32'b00000000000000000000000000000000;
		mem_arr[31]=32'b00000000000000000000000000000000;
	end
	 
    // initial begin
    //     $readmemh("file.txt", mem_arr);
    // end

    always @(MemRW) begin
        if (MemRW==read) begin
            dataB=mem_arr[addr[31:2]];
        end else begin
            dataB = 32'h00000000;
        end
    end

    always @(posedge clk) begin
        if (MemRW==write) begin
            mem_arr[addr[31:2]]<=dataW;
            //$memwriteh("file.txt", mem_arr);
        end
    end
endmodule